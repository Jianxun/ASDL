* SPICE netlist generated from ASDL
* Design: None
* Top module: inverter
* Author: None
* Date: None
* Revision: None

* Hierarchical module subcircuit definitions
* .subckt inverter in out vdd vss
  m1 out in vss vss nmos L=0.18u W=1u
  m2 out in vdd vdd pmos L=0.18u W=2u
* .ends


.end