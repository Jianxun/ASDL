Xdut IREF IOUT_P IOUT_N VSS current_mirror_array

* GF180MCU Model Card:
.include PDK_MODEL_PATH/design.ngspice
.lib PDK_MODEL_PATH/sm141064.ngspice typical

X_MN1 VSS VSS VSS VSS nfet_03v3 L=0.2u W=5u NF=2 m=1
* ===============================================
* current_mirror_array
.subckt current_mirror_array IREF IOUT_P IOUT_N VSS

X_MN_REF IREF IREF VSS VSS nfet_03v3 L=0.2u W=5u NF=2 m=1
X_MN_OUT_P IOUT_P IREF VSS VSS nfet_03v3 L=0.2u W=5u NF=1 m=1
X_MN_OUT_N IOUT_N IREF VSS VSS nfet_03v3 L=0.2u W=5u NF=1 m=1
.ends current_mirror_array

.end