
    * ---------------- Model Files ----------------
    .include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
    .lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
    
    * ---------------- Power Supplies ----------------
    V_vss vss 0 0
    V_vdd vdd 0 3.3
    
    * ---------------- Single Pulse Stimulus ----------------
    V_in in 0 PULSE(0 3.3 2e-09 5e-11 5e-11 1e-08 1)
    
    * ---------------- Transient Analysis ----------------
    .control
    save all
    TRAN 1e-11 2e-08 0
    write /foss/designs/simulations/inverter_asdl/test_prop_delay/prop_delay.raw
    .endc

    * SPICE netlist generated from ASDL
* Design: Basic CMOS inverter
* Top module: inverter
* Author: ASDL
* Date: 2024-03-19
* Revision: v0.4

* Model subcircuit definitions
* NMOS transistor unit cell
.subckt nmos_unit G D S B
  .param M=1
  .param nf=2
  .param L=0.5u
  .param W=4u
  MN D G S B nfet_03v3 L={L} W={W} nf={nf} M={M} ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0
.ends

* PMOS transistor unit cell
.subckt pmos_unit G D S B
  .param M=1
  .param nf=2
  .param L=0.5u
  .param W=5u
  MP D G S B pfet_03v3 L={L} W={W} nf={nf} M={M} ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0
.ends

* Basic CMOS inverter with PMOS pull-up and NMOS pull-down
.subckt inverter in out vss vdd
  .param M=1
  X_MP in out vdd vdd pmos_unit M=2
  X_MN in out vss vss nmos_unit M=2
.ends

* Main circuit instantiation
XMAIN in out vss vdd inverter

.end