* SPICE netlist generated from ASDL
* Design: Two-stage Miller-compensated operational transconductance amplifier
* Top module: two_stage_ota
* Author: ASDL
* Date: 2025-06-14
* Revision: v0.4

* Model subcircuit definitions
* Small resistor net jumper
.subckt jumper plus minus
  R1 plus minus R=100m
.ends

* NMOS transistor unit cell
.subckt nmos_unit G D S B
  .param M=1
  MN D G S B nfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* PMOS transistor unit cell
.subckt pmos_unit G D S B
  .param M=1
  MP D G S B pfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* Miller compensation capacitor
.subckt comp_cap plus minus
  C1 plus minus C=1p
.ends

* Miller compensation resistor
.subckt comp_res plus minus
  R1 plus minus R=1k
.ends

* Bias generator
.subckt bias_gen ibias vbn vss vdd
  X_MN_BIAS vbn vbn vss vss nmos_unit M=1
  X_J1 ibias vbn jumper
.ends

* 5-transistor OTA: differential pair with current mirror load
.subckt ota_5t in_p in_n out vbn vss vdd
  .param M=2
  * NMOS input transistors
  X_MN_P in_p vd tail vss nmos_unit M={M}
  * NMOS input transistors
  X_MN_N in_n out tail vss nmos_unit M={M}
  * NMOS tail current source
  X_MN_TAIL vbn tail vss vss nmos_unit M={M}*2
  * PMOS current mirror load
  X_MP_P vd vd vdd vdd pmos_unit M={M}*3
  * PMOS current mirror load
  X_MP_N vd out vdd vdd pmos_unit M={M}*3
.ends

* Second stage: PMOS Common source amplifier with NMOS current source load
.subckt common_source_pmos in out vbn vss vdd
  .param M=4
  X_MP_CS in out vdd vdd pmos_unit M={M}*3
  X_MN_LOAD vbn out vss vss nmos_unit M={M}
.ends

* Miller compensation network
.subckt miller_comp plus minus
  X_CC plus v_int comp_cap
  X_RC v_int minus comp_res
.ends

* Two-stage Miller-compensated operational transconductance amplifier
.subckt two_stage_ota in_p in_n out ibias vss vdd
  .param M_first_stage=2
  .param M_second_stage=4
  X_BIAS_GEN ibias vbn vss vdd bias_gen
  X_FIRST_STAGE in_n in_p first_stage_out vbn vss vdd ota_5t M={M_first_stage}
  X_SECOND_STAGE first_stage_out out vbn vss vdd common_source_pmos M={M_second_stage}
  X_COMP first_stage_out out miller_comp
.ends

* Main circuit instantiation
XMAIN in_p in_n out ibias vss vdd two_stage_ota

.end