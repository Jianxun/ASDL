* SPICE netlist generated from ASDL
* Design: A collection of differential pairs
* Top module: diff_pair
* Author: ASDL
* Date: 2025-06-25
* Revision: v0.1

* Model subcircuit definitions
* NMOS transistor unit cell
.subckt nmos_unit G D S B
  .param M=1
  MN D G S B nfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0
.ends

* PMOS transistor unit cell
.subckt pmos_unit G D S B
  .param M=1
  MP D G S B pfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0
.ends

* Miller compensation capacitor
.subckt cap plus minus
  C1 plus minus C=1p
.ends

* Miller compensation resistor
.subckt res plus minus
  R1 plus minus R=1k
.ends

* Differential pair NMOS
.subckt diff_pair_nmos vdd inp inn outp outn vbn vss
  .param R=1k
  .param M=1
  X_MN_DPP inp outn tail vss nmos_unit M={M}
  X_MN_DPN inn outp tail vss nmos_unit M={M}
  X_M_TAIL vbn tail vss vss nmos_unit M={M}
  X_R_LOADP vdd outn res R={R}
  X_R_LOADN vdd outp res R={R}
.ends


.end