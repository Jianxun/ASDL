* ===============================================
subckt tb

M_MN1 d g s b nfet_03v3 L=0.5u W=5u NF=2 m=1
R_R1 g s 1k





ends