* SPICE netlist generated from ASDL
* Design: Demonstration of unified ASDL architecture with primitive and hierarchical modules
* Top module: two_stage_buffer
* Author: ASDL Unified Architecture Demo
* Date: 2024-03-15
* Revision: 1.0

* PDK model includes
.include "gf180mcu_fd_pr/models/ngspice/design.ngspice"

* Hierarchical module subcircuit definitions
* CMOS inverter using PDK primitives
.subckt inverter in out vdd vss
  XMN out in vss vss nfet_03v3 L=0.28u W=3u m=1
  XMP out in vdd vdd pfet_03v3 L=0.28u W=6u m=2
.ends

* RC filter configured for buffer application
.subckt buffer_rc_filter in out gnd
  RR1 in out 5k TC1=0 TC2=0
  CC1 out gnd 50p
.ends

* NMOS current mirror with 1:2:4 current ratios
.subckt current_mirror iref iout1 iout2 vss
  XM_REF iref iref vss vss nfet_03v3 L=0.28u W=3u m=1
  XM_OUT1 iout1 iref vss vss nfet_03v3 L=0.28u W=3u m=2
  XM_OUT2 iout2 iref vss vss nfet_03v3 L=0.28u W=3u m=4
.ends

* Two-stage buffer with RC filter - demonstrates mixed hierarchy
.subckt two_stage_buffer in out vdd vss
  X_INV1 in stage1_out vdd vss inverter
  X_FILTER stage1_out filtered_out vss buffer_rc_filter
  * First parallel inverter for drive strength
  X_INV2A filtered_out out vdd vss inverter
  * Second parallel inverter for drive strength
  X_INV2B filtered_out out vdd vss inverter
  * Demonstration current mirror - would connect to bias circuitry
  X_CM1 vss vss vss vss current_mirror
.ends

* Main circuit instantiation
XMAIN in out vdd vss two_stage_buffer

.end