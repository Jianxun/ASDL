🎉 Successfully generated: examples/two_stage_ota.spice
