
    * ---------------- Model Files ----------------
    .include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
    .lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
    
    * ---------------- Power Supplies ----------------
    V_vss vss 0 0
    V_vdd vdd 0 3.3
    
    * ---------------- DC Sweep Stimulus ----------------
    V_in in 0 0
    
    * ---------------- DC Sweep Analysis ----------------
    .control
    save all
    DC V_in 0 3.3 0.01
    write /foss/designs/simulations/inverter_asdl/test_dc_transfer/dc_transfer.raw
    .endc

    * SPICE netlist generated from ASDL
* Design: Basic CMOS inverter
* Top module: inverter
* Author: ASDL
* Date: 2024-03-19
* Revision: v0.4

* Model subcircuit definitions
* NMOS transistor unit cell
.subckt nmos_unit G D S B
  .param M=1
  MN D G S B nfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* PMOS transistor unit cell
.subckt pmos_unit G D S B
  .param M=1
  MP D G S B pfet_03v3 L=0.5u W=5u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* Basic CMOS inverter with PMOS pull-up and NMOS pull-down
.subckt inverter in out vss vdd
  .param M=1
  X_MP in out vdd vdd pmos_unit M=2
  X_MN in out vss vss nmos_unit M=2
.ends

* Main circuit instantiation
XMAIN in out vss vdd inverter

.end