* SPICE netlist generated from ASDL
* Design: NMOS differential pair with resistor loads - Pattern expansion test circuit
* Author: ASDL Test Suite
* Date: 2024-03-19
* Revision: v0.4

* Model subcircuit definitions
* NMOS transistor unit cell
.subckt nmos_unit G D S B
  .param M=1
  MN D G S B nfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* Resistor unit cell
.subckt resistor_unit plus minus
  .param R=10k
  R1 plus minus ppolyf_u L=2u W=1u m=1 R={R}
.ends

* NMOS differential pair with resistor loads demonstrating pattern expansion
.subckt diff_pair_nmos in_n in_p iref out_n out_p tail vdd vss
  X_MN_P in_p out_p tail vss nmos_unit M=$M_diff
  X_MN_N in_p out_p tail vss nmos_unit M=$M_diff
  X_RL_P vdd out_p resistor_unit R=$R_load
  X_RL_N vdd out_p resistor_unit R=$R_load
  X_M_DIODE bias_gate bias_gate vss vss nmos_unit M=$M_diode
  X_M_MIRROR bias_gate tail vss vss nmos_unit M=$M_mirror
.ends

* Main circuit instantiation
XMAIN in_n in_p iref out_n out_p tail vdd vss diff_pair_nmos

.end