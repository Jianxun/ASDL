* SPICE netlist generated from ASDL
* Design: Gray & Meyer 6th edition
Fig. 3.12
Resistive load common-source amplifier

* Top module: cs_amplifier
* Author: None
* Date: None
* Revision: None

* Hierarchical module subcircuit definitions
* Resistive load common-source amplifier
* .subckt cs_amplifier vdd vss vin vout
  X_mn1 vout vin vss vss nfet_03v3 L=0.28u W=3u nf=2 m=1
+ ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' 
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' 
+ nrd='0.18u / W' nrs='0.18u / W' 
+ sa=0 sb=0 sd=0

  rd vdd vout 10k

* .ends


.end