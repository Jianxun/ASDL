* SPICE netlist generated from ASDL
* Design: Two-stage Miller-compensated operational transconductance amplifier
* Author: ASDL
* Date: 2025-06-14
* Revision: v0.4

* Model subcircuit definitions
* Small resistor net jumper
.subckt jumper plus minus
  R1 plus minus R=100m
.ends

* NMOS transistor unit cell
.subckt nmos_unit G D S B
  .param M=1
  MN D G S B nfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* PMOS transistor unit cell
.subckt pmos_unit G D S B
  .param M=1
  MP D G S B pfet_03v3 L=0.5u W=4u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 M={M}
.ends

* Miller compensation capacitor
.subckt comp_cap plus minus
  C1 plus minus C=1p
.ends

* Miller compensation resistor
.subckt comp_res plus minus
  R1 plus minus R=1k
.ends

* Bias generator
.subckt bias_gen ibias vbn vdd vss
  X_MN_BIAS vbn vbn vss vss nmos_unit M=1
  X_J1 ibias vbn jumper
.ends

* 5-transistor OTA: differential pair with current mirror load
.subckt ota_5t in_n in_p out vbn vdd vss
  .param M=2
  * NMOS input transistors
  X_MN_P in_p vd tail vss nmos_unit M={M}
  * NMOS input transistors
  X_MN_N in_p vd tail vss nmos_unit M={M}
  * NMOS tail current source
  X_MN_TAIL vbn tail vss vss nmos_unit M={M}*2
  * PMOS current mirror load
  X_MP_P out_n out_p vdd vdd pmos_unit M={M}*3
  * PMOS current mirror load
  X_MP_N out_n out_p vdd vdd pmos_unit M={M}*3
.ends

* Second stage: PMOS Common source amplifier with NMOS current source load
.subckt common_source_pmos in out vbn vdd vss
  .param M=4
  X_MP_CS in out vdd vdd pmos_unit M={M}*3
  X_MN_LOAD vbn out vss vss nmos_unit M={M}
.ends

* Miller compensation network
.subckt miller_comp minus plus
  X_CC plus v_int comp_cap
  X_RC v_int minus comp_res
.ends

* Two-stage Miller-compensated operational transconductance amplifier
.subckt two_stage_ota ibias in_n in_p out vdd vss
  .param M.first_stage=2
  .param M.second_stage=4
  X_FIRST_STAGE in_p in_n first_stage_out vbn vdd vss ota_5t
  X_SECOND_STAGE first_stage_out out vbn vdd vss common_source_pmos
  X_COMP UNCONNECTED UNCONNECTED miller_comp
.ends

* Main circuit instantiation
XMAIN ibias in_n in_p out vdd vss two_stage_ota

.end