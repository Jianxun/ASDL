* SPICE netlist generated from ASDL
* Design: Basic CMOS inverter
* Top module: inverter
* Author: ASDL
* Date: 2024-03-19
* Revision: v0.4

* Hierarchical module subcircuit definitions
* Basic CMOS inverter with PMOS pull-up and NMOS pull-down
.subckt inverter 
* ERROR G0401: unknown model 'pmos_unit'
* ERROR G0401: unknown model 'nmos_unit'
.ends


.end