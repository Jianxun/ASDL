* SPICE netlist generated from ASDL
* Design: Test ASDL file
* Top module: test
* Author: None
* Date: None
* Revision: None

* Hierarchical module subcircuit definitions
* .subckt test in out
  vgs g vss DC 1

  vds d vss DC 0.5

  vss vss GND DC 0.0

  X_m1 d g vss vss nfet_03v3 L=0.28u W=3u nf=2 m=1
+ ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' 
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' 
+ nrd='0.18u / W' nrs='0.18u / W' 
+ sa=0 sb=0 sd=0

  .include ./gf180mcu/ngspice/design.ngspice
.lib ./gf180mcu/ngspice/sm141064.ngspice typical

  .control
save all
dc vds 0 3.3 0.05
*write to raw file
write sim_dc_results.raw
.endc
* .ends


.end